module tb();
int a;
intial begin
 a=10;
 end
 $monitor(a);
 endmodule
